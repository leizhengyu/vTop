// =====HEAD BEGIN ===============
// FileName  : aasdf
// Author    : liuzhiyong
// BuildTime : 2015-3-15
// =====HEAD END =================

module MODULE
(
// =====PORTS BEGIN ==============
// =====PORTS END ================
);
// =====WIRES BEGIN ==============
// =====WIRES END ================

// =====USERDEFINED BEGIN ========
// =====USERDEFINED END ==========

// =====INSTANCES BEGIN ==========
// =====INSTANCES END ============

// =====DEFINES BEGIN ============
// =====DEFINES END ==============

// =====UI BEGIN =================
// =====UI END ===================

endmodule
